library ieee;
use ieee.std_logic_1164.all;

entity thunderbird_fsm is
	port(
		i_clk, i_reset 	: in std_logic;  
		i_left, i_right 	: in std_logic; 
		o_lights_L 			: out std_logic_vector(2 downto 0); -- leds
		o_lights_R 			: out std_logic_vector(2 downto 0) -- leds
		);
end thunderbird_fsm;

architecture behaviour of thunderbird_fsm is
	
	type lights_state is (OFF, Flash, R1, R2, R3, L1, L2, L3);
   signal next_state, current_state : lights_state;

	begin
 
	-- current state logic defined below
	process (i_clk, i_reset)
		begin
		
			if(i_reset = '1') then
				current_state <= OFF;
			elsif rising_edge(i_clk) then
				current_state <= next_state;
			end if;
			
		end process;
	
	-- next state logic defined below
	process(current_state, i_left, i_right)
		begin
		case current_state is
			when OFF => if ((i_left = '1') and (i_right = '0')) then next_state <= L1;
							elsif ((i_left = '0') and (i_right = '1'))  then next_state <= R1;
							elsif((i_left = '1') and (i_right = '1'))  then next_state <= Flash;
							else next_state <= OFF;
							end if;
							
			when R1 => next_state <= R2;										
			
			when R2 => next_state <= R3;
							
			when R3 => next_state <= OFF;
							
			when L1 => next_state <= L2;
							
			when L2 => next_state <= L3;
							
			when L3 => next_state <= OFF;
							
			when Flash => next_state <= OFF;
							
			when others => next_state <= OFF;
			
		end case;
	end process;

	-- Output logic defined below
	
	o_lights_R <= "100" when (current_state = R1) else
					  "110" when (current_state = R2) else
					  "111" when ((current_state = R3) or (current_state = Flash)) else
					  "000" when (current_state = OFF);
	
	o_lights_L <= "001" when (current_state = L1) else
					  "011" when (current_state = L2) else
					  "111" when ((current_state = L3) or (current_state = Flash)) else
					  "000" when (current_state = OFF);
	
						
	
end behaviour;